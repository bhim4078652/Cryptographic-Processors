module decryptRound(i_clk,i_rst,in,i_key,out);
input i_clk,i_rst;
input [127:0] in;
output [127:0] out;
input [127:0] i_key;
wire [127:0] w_afterSubBytes;
wire [127:0] w_afterShiftRows;
wire [127:0] w_afterAddroundi_key;

inverseShiftRows r(in,w_afterShiftRows);
inverseSubBytes s(w_afterShiftRows,w_afterSubBytes);
addRoundKey b(i_clk,i_rst,w_afterSubBytes,w_afterAddroundi_key,i_key);
inverseMixColumns m(w_afterAddroundi_key,out);
		
endmodule